module notGate(x,y);
	input x;
	output y;
	assign y = ~x;
endmodule
